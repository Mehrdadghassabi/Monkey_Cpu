
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

entity Rom is
port (
 pc: in std_logic_vector(15 downto 0);
 result   : in  STD_LOGIC_VECTOR(15 downto 0);
 datins: out  std_logic_vector(31 downto 0)
);
end Rom;

architecture Behavioral of Rom is
 type ROM_type is array (0 to 63 ) of std_logic_vector(31 downto 0);
 type RAM_type is array (0 to 15 ) of std_logic_vector(15 downto 0);
 constant rom_ins: ROM_type:=(
   "11111111111111110000000011110011",
   "11111111100000000000000011011111",
   "11111111111111111111111110000110",
   "11111111111111111111111101111100",
   "11111111101000000000000011110011",
   "11111111100000000000000011011111",
   "11111111111111111111111110000110",
   "11111111111111111111111101111100",
   "11111111001001100000000011110011",
   "11111111100000000000000011011111",
   "11111111111111111111111110000110",
   "11111111111111111111111101111100",
   "11111111000000000000000011110011",
   "11111111011101000000000011011111",
   "11111111111111111111111110000110",
   "11111111111111111111111101111100",
   "11111111000000000000000011110011",
   "11111111000100110000000011011111",
   "11111111111111111111111110000110",
   "11111111111111111111111101111100",
   "11111111001001100000000011110011",
   "11111111111111111111111111011111",
   "11111111111111111111111110000110",
   "11111111111111111111111101111100",
   "11111111111111111111111111110011",
   "11111111001011010000000011011111",
   "11111111111111111111111110000110",
   "11111111111111111111111101111100",
   "11111111111111111111111111110011",
   "11111111001101001000000011011111",
   "11111111111111111111111110000110",
   "11111111111111111111111101111100",
   "11111111000000000000000011110011",
   "11111111000000000000000011011111",
   "11111111111111111111111110000110",
   "11111111111111111111111101111100",
   "11111111111111111111111100001101",
   "00000000000000000000000000000000",	
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
	"00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000"
  );
  signal ram_data: RAM_type:=(
   "0000000000000000",
   "0000000000000000",
   "0000000000000000",
	"0000000000000000",
   "0000000000000000",
   "0000000000000000",
	"0000000000000000",
   "0000000000000000",
   "0000000000000000",
	"0000000000000000",
   "0000000000000000",
   "0000000000000000",
	"0000000000000000",
   "0000000000000000",
   "0000000000000000",
	"0000000000000000"  
  );
begin
  
  datins <= rom_ins(to_integer(unsigned(pc)));
  ram_data(to_integer(unsigned(pc)))<= result ;

end Behavioral;


